module ALU(
  input  [3:0]  io_func, // @[common/src/main/scala/riscv/core/ALU.scala 27:14]
  input  [31:0] io_op1, // @[common/src/main/scala/riscv/core/ALU.scala 27:14]
  input  [31:0] io_op2, // @[common/src/main/scala/riscv/core/ALU.scala 27:14]
  output [31:0] io_result // @[common/src/main/scala/riscv/core/ALU.scala 27:14]
);
  wire [31:0] _io_result_T_1 = io_op1 + io_op2; // @[common/src/main/scala/riscv/core/ALU.scala 39:27]
  wire [31:0] _io_result_T_3 = io_op1 - io_op2; // @[common/src/main/scala/riscv/core/ALU.scala 42:27]
  wire [62:0] _GEN_10 = {{31'd0}, io_op1}; // @[common/src/main/scala/riscv/core/ALU.scala 45:27]
  wire [62:0] _io_result_T_5 = _GEN_10 << io_op2[4:0]; // @[common/src/main/scala/riscv/core/ALU.scala 45:27]
  wire [31:0] _io_result_T_6 = io_op1; // @[common/src/main/scala/riscv/core/ALU.scala 48:27]
  wire [31:0] _io_result_T_7 = io_op2; // @[common/src/main/scala/riscv/core/ALU.scala 48:43]
  wire [31:0] _io_result_T_9 = io_op1 ^ io_op2; // @[common/src/main/scala/riscv/core/ALU.scala 51:27]
  wire [31:0] _io_result_T_10 = io_op1 | io_op2; // @[common/src/main/scala/riscv/core/ALU.scala 54:27]
  wire [31:0] _io_result_T_11 = io_op1 & io_op2; // @[common/src/main/scala/riscv/core/ALU.scala 57:27]
  wire [31:0] _io_result_T_13 = io_op1 >> io_op2[4:0]; // @[common/src/main/scala/riscv/core/ALU.scala 60:27]
  wire [31:0] _io_result_T_17 = $signed(io_op1) >>> io_op2[4:0]; // @[common/src/main/scala/riscv/core/ALU.scala 63:52]
  wire  _GEN_0 = 4'ha == io_func & io_op1 < io_op2; // @[common/src/main/scala/riscv/core/ALU.scala 36:13 37:19 66:17]
  wire [31:0] _GEN_1 = 4'h9 == io_func ? _io_result_T_17 : {{31'd0}, _GEN_0}; // @[common/src/main/scala/riscv/core/ALU.scala 37:19 63:17]
  wire [31:0] _GEN_2 = 4'h8 == io_func ? _io_result_T_13 : _GEN_1; // @[common/src/main/scala/riscv/core/ALU.scala 37:19 60:17]
  wire [31:0] _GEN_3 = 4'h7 == io_func ? _io_result_T_11 : _GEN_2; // @[common/src/main/scala/riscv/core/ALU.scala 37:19 57:17]
  wire [31:0] _GEN_4 = 4'h6 == io_func ? _io_result_T_10 : _GEN_3; // @[common/src/main/scala/riscv/core/ALU.scala 37:19 54:17]
  wire [31:0] _GEN_5 = 4'h5 == io_func ? _io_result_T_9 : _GEN_4; // @[common/src/main/scala/riscv/core/ALU.scala 37:19 51:17]
  wire [31:0] _GEN_6 = 4'h4 == io_func ? {{31'd0}, $signed(_io_result_T_6) < $signed(_io_result_T_7)} : _GEN_5; // @[common/src/main/scala/riscv/core/ALU.scala 37:19 48:17]
  wire [62:0] _GEN_7 = 4'h3 == io_func ? _io_result_T_5 : {{31'd0}, _GEN_6}; // @[common/src/main/scala/riscv/core/ALU.scala 37:19 45:17]
  wire [62:0] _GEN_8 = 4'h2 == io_func ? {{31'd0}, _io_result_T_3} : _GEN_7; // @[common/src/main/scala/riscv/core/ALU.scala 37:19 42:17]
  wire [62:0] _GEN_9 = 4'h1 == io_func ? {{31'd0}, _io_result_T_1} : _GEN_8; // @[common/src/main/scala/riscv/core/ALU.scala 37:19 39:17]
  assign io_result = _GEN_9[31:0];
endmodule
module ALUControl(
  input  [6:0] io_opcode, // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 21:14]
  input  [2:0] io_funct3, // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 21:14]
  input  [6:0] io_funct7, // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 21:14]
  output [3:0] io_alu_funct // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 21:14]
);
  wire [3:0] _io_alu_funct_T_1 = io_funct7[5] ? 4'h9 : 4'h8; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 66:41]
  wire  _io_alu_funct_T_2 = 3'h1 == io_funct3; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire [1:0] _io_alu_funct_T_3 = 3'h1 == io_funct3 ? 2'h3 : 2'h1; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire  _io_alu_funct_T_4 = 3'h2 == io_funct3; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire [2:0] _io_alu_funct_T_5 = 3'h2 == io_funct3 ? 3'h4 : {{1'd0}, _io_alu_funct_T_3}; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire  _io_alu_funct_T_6 = 3'h3 == io_funct3; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire [3:0] _io_alu_funct_T_7 = 3'h3 == io_funct3 ? 4'ha : {{1'd0}, _io_alu_funct_T_5}; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire  _io_alu_funct_T_8 = 3'h4 == io_funct3; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire [3:0] _io_alu_funct_T_9 = 3'h4 == io_funct3 ? 4'h5 : _io_alu_funct_T_7; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire  _io_alu_funct_T_10 = 3'h6 == io_funct3; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire [3:0] _io_alu_funct_T_11 = 3'h6 == io_funct3 ? 4'h6 : _io_alu_funct_T_9; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire  _io_alu_funct_T_12 = 3'h7 == io_funct3; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire [3:0] _io_alu_funct_T_13 = 3'h7 == io_funct3 ? 4'h7 : _io_alu_funct_T_11; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire  _io_alu_funct_T_14 = 3'h5 == io_funct3; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire [3:0] _io_alu_funct_T_15 = 3'h5 == io_funct3 ? _io_alu_funct_T_1 : _io_alu_funct_T_13; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 48:62]
  wire [1:0] _io_alu_funct_T_17 = io_funct7[5] ? 2'h2 : 2'h1; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 83:43]
  wire [1:0] _io_alu_funct_T_21 = _io_alu_funct_T_2 ? 2'h3 : _io_alu_funct_T_17; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 77:62]
  wire [2:0] _io_alu_funct_T_23 = _io_alu_funct_T_4 ? 3'h4 : {{1'd0}, _io_alu_funct_T_21}; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 77:62]
  wire [3:0] _io_alu_funct_T_25 = _io_alu_funct_T_6 ? 4'ha : {{1'd0}, _io_alu_funct_T_23}; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 77:62]
  wire [3:0] _io_alu_funct_T_27 = _io_alu_funct_T_8 ? 4'h5 : _io_alu_funct_T_25; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 77:62]
  wire [3:0] _io_alu_funct_T_29 = _io_alu_funct_T_10 ? 4'h6 : _io_alu_funct_T_27; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 77:62]
  wire [3:0] _io_alu_funct_T_31 = _io_alu_funct_T_12 ? 4'h7 : _io_alu_funct_T_29; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 77:62]
  wire [3:0] _io_alu_funct_T_33 = _io_alu_funct_T_14 ? _io_alu_funct_T_1 : _io_alu_funct_T_31; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 77:62]
  wire [3:0] _GEN_0 = 7'h33 == io_opcode ? _io_alu_funct_T_33 : 4'h1; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 43:16 45:21 77:20]
  assign io_alu_funct = 7'h13 == io_opcode ? _io_alu_funct_T_15 : _GEN_0; // @[1-single-cycle/src/main/scala/riscv/core/ALUControl.scala 45:21 48:20]
endmodule
module Execute(
  input         clock,
  input         reset,
  input  [31:0] io_instruction, // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 45:14]
  input  [31:0] io_instruction_address, // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 45:14]
  input  [31:0] io_reg1_data, // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 45:14]
  input  [31:0] io_reg2_data, // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 45:14]
  input  [31:0] io_immediate, // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 45:14]
  input         io_aluop1_source, // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 45:14]
  input         io_aluop2_source, // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 45:14]
  output [31:0] io_mem_alu_result, // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 45:14]
  output        io_if_jump_flag, // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 45:14]
  output [31:0] io_if_jump_address // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 45:14]
);
  wire [3:0] alu_io_func; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 65:24]
  wire [31:0] alu_io_op1; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 65:24]
  wire [31:0] alu_io_op2; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 65:24]
  wire [31:0] alu_io_result; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 65:24]
  wire [6:0] alu_ctrl_io_opcode; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 66:24]
  wire [2:0] alu_ctrl_io_funct3; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 66:24]
  wire [6:0] alu_ctrl_io_funct7; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 66:24]
  wire [3:0] alu_ctrl_io_alu_funct; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 66:24]
  wire [6:0] opcode = io_instruction[6:0]; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 60:30]
  wire [2:0] funct3 = io_instruction[14:12]; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 61:30]
  wire  _branchCondition_T = io_reg1_data == io_reg2_data; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 96:47]
  wire  _branchCondition_T_1 = io_reg1_data != io_reg2_data; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 99:47]
  wire  _branchCondition_T_4 = $signed(io_reg1_data) < $signed(io_reg2_data); // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 103:54]
  wire  _branchCondition_T_7 = $signed(io_reg1_data) >= $signed(io_reg2_data); // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 106:54]
  wire  _branchCondition_T_8 = io_reg1_data < io_reg2_data; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 110:47]
  wire  _branchCondition_T_9 = io_reg1_data >= io_reg2_data; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 113:47]
  wire  _branchCondition_T_13 = 3'h1 == funct3 ? _branchCondition_T_1 : 3'h0 == funct3 & _branchCondition_T; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 90:51]
  wire  _branchCondition_T_15 = 3'h4 == funct3 ? _branchCondition_T_4 : _branchCondition_T_13; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 90:51]
  wire  _branchCondition_T_17 = 3'h5 == funct3 ? _branchCondition_T_7 : _branchCondition_T_15; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 90:51]
  wire  _branchCondition_T_19 = 3'h6 == funct3 ? _branchCondition_T_8 : _branchCondition_T_17; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 90:51]
  wire  branchCondition = 3'h7 == funct3 ? _branchCondition_T_9 : _branchCondition_T_19; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 90:51]
  wire  isBranch = opcode == 7'h63; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 116:25]
  wire  isJal = opcode == 7'h6f; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 117:25]
  wire  isJalr = opcode == 7'h67; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 118:25]
  wire [31:0] branchTarget = io_instruction_address + io_immediate; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 131:45]
  wire [31:0] jalrSum = io_reg1_data + io_immediate; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 139:35]
  wire [31:0] jalrTarget = {jalrSum[31:1],1'h0}; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 143:23]
  wire  branchTaken = isBranch & branchCondition; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 145:30]
  ALU alu ( // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 65:24]
    .io_func(alu_io_func),
    .io_op1(alu_io_op1),
    .io_op2(alu_io_op2),
    .io_result(alu_io_result)
  );
  ALUControl alu_ctrl ( // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 66:24]
    .io_opcode(alu_ctrl_io_opcode),
    .io_funct3(alu_ctrl_io_funct3),
    .io_funct7(alu_ctrl_io_funct7),
    .io_alu_funct(alu_ctrl_io_alu_funct)
  );
  assign io_mem_alu_result = alu_io_result; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 79:21]
  assign io_if_jump_flag = branchTaken | isJal | isJalr; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 146:43]
  assign io_if_jump_address = isJalr ? jalrTarget : branchTarget; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 147:28]
  assign alu_io_func = alu_ctrl_io_alu_funct; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 73:15]
  assign alu_io_op1 = io_aluop1_source ? io_instruction_address : io_reg1_data; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 74:19]
  assign alu_io_op2 = io_aluop2_source ? io_immediate : io_reg2_data; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 75:19]
  assign alu_ctrl_io_opcode = io_instruction[6:0]; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 60:30]
  assign alu_ctrl_io_funct3 = io_instruction[14:12]; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 61:30]
  assign alu_ctrl_io_funct7 = io_instruction[31:25]; // @[1-single-cycle/src/main/scala/riscv/core/Execute.scala 62:30]
endmodule
