module InstructionDecode(
  input         clock,
  input         reset,
  input  [31:0] io_instruction, // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 150:14]
  output [4:0]  io_regs_reg1_read_address, // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 150:14]
  output [4:0]  io_regs_reg2_read_address, // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 150:14]
  output [31:0] io_ex_immediate, // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 150:14]
  output        io_ex_aluop1_source, // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 150:14]
  output        io_ex_aluop2_source, // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 150:14]
  output        io_memory_read_enable, // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 150:14]
  output        io_memory_write_enable, // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 150:14]
  output [1:0]  io_wb_reg_write_source, // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 150:14]
  output        io_reg_write_enable, // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 150:14]
  output [4:0]  io_reg_write_address // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 150:14]
);
  wire [6:0] opcode = io_instruction[6:0]; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 166:32]
  wire [4:0] rs1 = io_instruction[19:15]; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 167:32]
  wire [4:0] rs2 = io_instruction[24:20]; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 168:32]
  wire [4:0] rd = io_instruction[11:7]; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 169:32]
  wire  isLoad = opcode == 7'h3; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 171:25]
  wire  isStore = opcode == 7'h23; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 172:25]
  wire  isOpImm = opcode == 7'h13; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 173:25]
  wire  isOp = opcode == 7'h33; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 174:25]
  wire  isLui = opcode == 7'h37; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 175:25]
  wire  isAuipc = opcode == 7'h17; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 176:25]
  wire  isJal = opcode == 7'h6f; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 177:25]
  wire  isJalr = opcode == 7'h67; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 178:25]
  wire  isBranch = opcode == 7'h63; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 179:25]
  wire  _usesRs1_T_1 = isLoad | isStore | isOpImm; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 180:36]
  wire  usesRs1 = isLoad | isStore | isOpImm | isOp | isBranch | isJalr; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 180:67]
  wire  usesRs2 = isStore | isOp | isBranch; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 181:34]
  wire  _regWrite_T = isLoad | isOpImm; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 182:25]
  wire [1:0] _GEN_0 = isJal | isJalr ? 2'h2 : 2'h0; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 204:30 205:14 198:29]
  wire  _T_4 = _regWrite_T | isJalr; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 231:26]
  wire [1:0] _GEN_5 = isStore ? 2'h2 : {{1'd0}, _T_4}; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 234:17 235:13]
  wire [1:0] _GEN_6 = isBranch ? 2'h3 : _GEN_5; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 237:18 238:13]
  wire [2:0] _GEN_7 = isLui | isAuipc ? 3'h4 : {{1'd0}, _GEN_6}; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 240:26 241:13]
  wire [2:0] immKind = isJal ? 3'h5 : _GEN_7; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 243:15 244:13]
  wire [19:0] _immI_T_1 = io_instruction[31] ? 20'hfffff : 20'h0; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 269:9]
  wire [31:0] immI = {_immI_T_1,io_instruction[31:20]}; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 268:17]
  wire [31:0] immS = {_immI_T_1,io_instruction[31:25],rd}; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 279:17]
  wire [18:0] _immB_T_1 = io_instruction[31] ? 19'h7ffff : 19'h0; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 293:9]
  wire [31:0] immB = {_immB_T_1,io_instruction[31],io_instruction[7],io_instruction[30:25],io_instruction[11:8],1'h0}; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 292:17]
  wire [31:0] immU = {io_instruction[31:12],12'h0}; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 305:17]
  wire [10:0] _immJ_T_1 = io_instruction[31] ? 11'h7ff : 11'h0; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 315:9]
  wire [31:0] immJ = {_immJ_T_1,io_instruction[31],io_instruction[19:12],io_instruction[20],io_instruction[30:21],1'h0}; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 314:17]
  wire [31:0] _immediate_T_7 = 3'h1 == immKind ? immI : 32'h0; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 323:72]
  wire [31:0] _immediate_T_9 = 3'h2 == immKind ? immS : _immediate_T_7; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 323:72]
  wire [31:0] _immediate_T_11 = 3'h3 == immKind ? immB : _immediate_T_9; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 323:72]
  wire [31:0] _immediate_T_13 = 3'h4 == immKind ? immU : _immediate_T_11; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 323:72]
  assign io_regs_reg1_read_address = usesRs1 ? rs1 : 5'h0; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 247:35]
  assign io_regs_reg2_read_address = usesRs2 ? rs2 : 5'h0; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 248:35]
  assign io_ex_immediate = 3'h5 == immKind ? immJ : _immediate_T_13; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 323:72]
  assign io_ex_aluop1_source = isBranch | isAuipc | isJal; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 215:28]
  assign io_ex_aluop2_source = _usesRs1_T_1 | isBranch | isLui | isAuipc | isJal | isJalr; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 222:94]
  assign io_memory_read_enable = opcode == 7'h3; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 171:25]
  assign io_memory_write_enable = opcode == 7'h23; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 172:25]
  assign io_wb_reg_write_source = isLoad ? 2'h1 : _GEN_0; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 200:16 201:14]
  assign io_reg_write_enable = isLoad | isOpImm | isOp | isLui | isAuipc | isJal | isJalr; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 182:73]
  assign io_reg_write_address = io_instruction[11:7]; // @[1-single-cycle/src/main/scala/riscv/core/InstructionDecode.scala 169:32]
endmodule
